16 uid=11645753
26 mtime=1692274927.68242
27 atime=1692274927.681447
26 ctime=1692274927.68242
